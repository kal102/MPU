// qsys_top_mpu_ss_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module qsys_top_mpu_ss_0 (
		input  wire        clk_clk,                              //                    clk.clk
		input  wire        receive_startofpacket,                //                receive.startofpacket
		input  wire        receive_valid,                        //                       .valid
		output wire        receive_ready,                        //                       .ready
		input  wire [5:0]  receive_error,                        //                       .error
		input  wire [7:0]  receive_data,                         //                       .data
		input  wire        receive_endofpacket,                  //                       .endofpacket
		input  wire [1:0]  receive_empty,                        //                       .empty
		input  wire        reset_reset_n,                        //                  reset.reset_n
		input  wire        rx_mac_misc_connection_ff_rx_dsav,    // rx_mac_misc_connection.ff_rx_dsav
		input  wire        rx_mac_misc_connection_ff_rx_a_empty, //                       .ff_rx_a_empty
		input  wire        rx_mac_misc_connection_ff_rx_a_full,  //                       .ff_rx_a_full
		input  wire [17:0] rx_mac_misc_connection_rx_err_stat,   //                       .rx_err_stat
		input  wire [3:0]  rx_mac_misc_connection_rx_frm_type,   //                       .rx_frm_type
		output wire [31:0] transmit_data,                        //               transmit.data
		output wire        transmit_endofpacket,                 //                       .endofpacket
		output wire        transmit_error,                       //                       .error
		input  wire        transmit_ready,                       //                       .ready
		output wire        transmit_startofpacket,               //                       .startofpacket
		output wire        transmit_valid,                       //                       .valid
		output wire [1:0]  transmit_empty,                       //                       .empty
		output wire        tx_mac_misc_connection_ff_tx_crc_fwd, // tx_mac_misc_connection.ff_tx_crc_fwd
		input  wire        tx_mac_misc_connection_ff_tx_septy,   //                       .ff_tx_septy
		input  wire        tx_mac_misc_connection_ff_tx_uflow,   //                       .ff_tx_uflow
		input  wire        tx_mac_misc_connection_ff_tx_a_full,  //                       .ff_tx_a_full
		input  wire        tx_mac_misc_connection_ff_tx_a_empty  //                       .ff_tx_a_empty
	);

	wire         eth_rx_0_mpu_rx_buffer_a_b;     // eth_rx_0:buffer_a_b -> mpu_0:buffer_a_b
	wire         mpu_0_mpu_rx_mpu_ready;         // mpu_0:mpu_ready -> eth_rx_0:mpu_ready
	wire   [7:0] eth_rx_0_mpu_rx_buffer_a_data;  // eth_rx_0:buffer_a_data -> mpu_0:buffer_a_data
	wire   [4:0] eth_rx_0_mpu_rx_buffer_a_idx;   // eth_rx_0:buffer_a_idx -> mpu_0:buffer_a_idx
	wire   [7:0] eth_rx_0_mpu_rx_dim_y;          // eth_rx_0:dim_y -> mpu_0:dim_y_in
	wire   [7:0] eth_rx_0_mpu_rx_buffer_b_data;  // eth_rx_0:buffer_b_data -> mpu_0:buffer_b_data
	wire   [7:0] eth_rx_0_mpu_rx_dim_x;          // eth_rx_0:dim_x -> mpu_0:dim_x_in
	wire         eth_rx_0_mpu_rx_load;           // eth_rx_0:load -> mpu_0:load
	wire   [7:0] eth_rx_0_mpu_rx_pooling;        // eth_rx_0:pooling -> mpu_0:pooling
	wire  [23:0] eth_rx_0_mpu_rx_bias;           // eth_rx_0:bias -> mpu_0:bias
	wire   [4:0] eth_rx_0_mpu_rx_buffer_b_idx;   // eth_rx_0:buffer_b_idx -> mpu_0:buffer_b_idx
	wire         eth_rx_0_mpu_rx_buffer_ab_stop; // eth_rx_0:buffer_stop -> mpu_0:buffer_ab_stop
	wire   [7:0] eth_rx_0_mpu_rx_activation;     // eth_rx_0:activation -> mpu_0:activation
	wire         eth_rx_0_mpu_rx_multiply;       // eth_rx_0:multiply -> mpu_0:multiply
	wire   [7:0] mpu_0_mpu_tx_dim_y;             // mpu_0:dim_y_out -> eth_tx_0:dim_y
	wire   [7:0] mpu_0_mpu_tx_dim_x;             // mpu_0:dim_x_out -> eth_tx_0:dim_x
	wire         mpu_0_mpu_tx_data_available;    // mpu_0:data_available -> eth_tx_0:data_available
	wire         eth_tx_0_mpu_tx_buffer_c_stop;  // eth_tx_0:buffer_c_stop -> mpu_0:buffer_c_stop
	wire         mpu_0_mpu_tx_dim_error;         // mpu_0:dim_error -> eth_tx_0:dim_error
	wire         eth_tx_0_mpu_tx_tx_ready;       // eth_tx_0:tx_ready -> mpu_0:tx_ready
	wire  [23:0] mpu_0_mpu_tx_buffer_c_data;     // mpu_0:buffer_c_data -> eth_tx_0:buffer_c_data
	wire  [47:0] eth_rx_0_rx_tx_host_mac;        // eth_rx_0:host_mac -> eth_tx_0:host_mac
	wire   [7:0] eth_rx_0_rx_tx_rx_error;        // eth_rx_0:rx_error -> eth_tx_0:rx_error
	wire         rst_controller_reset_out_reset; // rst_controller:reset_out -> [eth_rx_0:rst_n, eth_tx_0:rst_n, mpu_0:rst_n]

	eth_rx #(
		.MMU_SIZE (10)
	) eth_rx_0 (
		.clk           (clk_clk),                              //                  clock.clk
		.rst_n         (~rst_controller_reset_out_reset),      //             reset_sink.reset_n
		.startofpacket (receive_startofpacket),                //                receive.startofpacket
		.valid         (receive_valid),                        //                       .valid
		.ready         (receive_ready),                        //                       .ready
		.error         (receive_error),                        //                       .error
		.data          (receive_data),                         //                       .data
		.endofpacket   (receive_endofpacket),                  //                       .endofpacket
		.mod           (receive_empty),                        //                       .empty
		.rx_error      (eth_rx_0_rx_tx_rx_error),              //                  rx_tx.rx_error
		.host_mac      (eth_rx_0_rx_tx_host_mac),              //                       .host_mac
		.dsav          (rx_mac_misc_connection_ff_rx_dsav),    // rx_mac_misc_connection.ff_rx_dsav
		.a_empty       (rx_mac_misc_connection_ff_rx_a_empty), //                       .ff_rx_a_empty
		.a_full        (rx_mac_misc_connection_ff_rx_a_full),  //                       .ff_rx_a_full
		.err_stat      (rx_mac_misc_connection_rx_err_stat),   //                       .rx_err_stat
		.frm_type      (rx_mac_misc_connection_rx_frm_type),   //                       .rx_frm_type
		.mpu_ready     (mpu_0_mpu_rx_mpu_ready),               //                 mpu_rx.mpu_ready
		.activation    (eth_rx_0_mpu_rx_activation),           //                       .activation
		.bias          (eth_rx_0_mpu_rx_bias),                 //                       .bias
		.buffer_a_b    (eth_rx_0_mpu_rx_buffer_a_b),           //                       .buffer_a_b
		.buffer_a_data (eth_rx_0_mpu_rx_buffer_a_data),        //                       .buffer_a_data
		.buffer_a_idx  (eth_rx_0_mpu_rx_buffer_a_idx),         //                       .buffer_a_idx
		.buffer_b_data (eth_rx_0_mpu_rx_buffer_b_data),        //                       .buffer_b_data
		.buffer_b_idx  (eth_rx_0_mpu_rx_buffer_b_idx),         //                       .buffer_b_idx
		.buffer_stop   (eth_rx_0_mpu_rx_buffer_ab_stop),       //                       .buffer_ab_stop
		.dim_x         (eth_rx_0_mpu_rx_dim_x),                //                       .dim_x
		.dim_y         (eth_rx_0_mpu_rx_dim_y),                //                       .dim_y
		.load          (eth_rx_0_mpu_rx_load),                 //                       .load
		.multiply      (eth_rx_0_mpu_rx_multiply),             //                       .multiply
		.pooling       (eth_rx_0_mpu_rx_pooling)               //                       .pooling
	);

	eth_tx eth_tx_0 (
		.rst_n          (~rst_controller_reset_out_reset),      //             reset_sink.reset_n
		.data           (transmit_data),                        //               transmit.data
		.endofpacket    (transmit_endofpacket),                 //                       .endofpacket
		.error          (transmit_error),                       //                       .error
		.ready          (transmit_ready),                       //                       .ready
		.startofpacket  (transmit_startofpacket),               //                       .startofpacket
		.wren           (transmit_valid),                       //                       .valid
		.mod            (transmit_empty),                       //                       .empty
		.host_mac       (eth_rx_0_rx_tx_host_mac),              //                  rx_tx.host_mac
		.rx_error       (eth_rx_0_rx_tx_rx_error),              //                       .rx_error
		.clk            (clk_clk),                              //                  clock.clk
		.crc_fwd        (tx_mac_misc_connection_ff_tx_crc_fwd), // tx_mac_misc_connection.ff_tx_crc_fwd
		.septy          (tx_mac_misc_connection_ff_tx_septy),   //                       .ff_tx_septy
		.uflow          (tx_mac_misc_connection_ff_tx_uflow),   //                       .ff_tx_uflow
		.a_full         (tx_mac_misc_connection_ff_tx_a_full),  //                       .ff_tx_a_full
		.a_empty        (tx_mac_misc_connection_ff_tx_a_empty), //                       .ff_tx_a_empty
		.buffer_c_data  (mpu_0_mpu_tx_buffer_c_data),           //                 mpu_tx.buffer_c_data
		.buffer_c_stop  (eth_tx_0_mpu_tx_buffer_c_stop),        //                       .buffer_c_stop
		.data_available (mpu_0_mpu_tx_data_available),          //                       .data_available
		.dim_error      (mpu_0_mpu_tx_dim_error),               //                       .dim_error
		.dim_x          (mpu_0_mpu_tx_dim_x),                   //                       .dim_x
		.dim_y          (mpu_0_mpu_tx_dim_y),                   //                       .dim_y
		.tx_ready       (eth_tx_0_mpu_tx_tx_ready)              //                       .tx_ready
	);

	mpu #(
		.VAR_SIZE  (8),
		.ACC_SIZE  (24),
		.MMU_SIZE  (10),
		.FIFO_SIZE (4)
	) mpu_0 (
		.clk            (clk_clk),                         //      clock.clk
		.rst_n          (~rst_controller_reset_out_reset), // reset_sink.reset_n
		.activation     (eth_rx_0_mpu_rx_activation),      //     mpu_rx.activation
		.bias           (eth_rx_0_mpu_rx_bias),            //           .bias
		.buffer_a_b     (eth_rx_0_mpu_rx_buffer_a_b),      //           .buffer_a_b
		.buffer_a_data  (eth_rx_0_mpu_rx_buffer_a_data),   //           .buffer_a_data
		.buffer_a_idx   (eth_rx_0_mpu_rx_buffer_a_idx),    //           .buffer_a_idx
		.buffer_ab_stop (eth_rx_0_mpu_rx_buffer_ab_stop),  //           .buffer_ab_stop
		.buffer_b_data  (eth_rx_0_mpu_rx_buffer_b_data),   //           .buffer_b_data
		.buffer_b_idx   (eth_rx_0_mpu_rx_buffer_b_idx),    //           .buffer_b_idx
		.dim_x_in       (eth_rx_0_mpu_rx_dim_x),           //           .dim_x
		.dim_y_in       (eth_rx_0_mpu_rx_dim_y),           //           .dim_y
		.load           (eth_rx_0_mpu_rx_load),            //           .load
		.multiply       (eth_rx_0_mpu_rx_multiply),        //           .multiply
		.pooling        (eth_rx_0_mpu_rx_pooling),         //           .pooling
		.mpu_ready      (mpu_0_mpu_rx_mpu_ready),          //           .mpu_ready
		.buffer_c_data  (mpu_0_mpu_tx_buffer_c_data),      //     mpu_tx.buffer_c_data
		.buffer_c_stop  (eth_tx_0_mpu_tx_buffer_c_stop),   //           .buffer_c_stop
		.data_available (mpu_0_mpu_tx_data_available),     //           .data_available
		.dim_error      (mpu_0_mpu_tx_dim_error),          //           .dim_error
		.dim_x_out      (mpu_0_mpu_tx_dim_x),              //           .dim_x
		.dim_y_out      (mpu_0_mpu_tx_dim_y),              //           .dim_y
		.tx_ready       (eth_tx_0_mpu_tx_tx_ready)         //           .tx_ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
